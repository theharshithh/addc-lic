module test_clt;            //test bench for the given QRS peak detection using CLT

  wire [31:0] out;          // the returned output is received in this array of wires
  reg [31:0] Yin;           // the input ECG value is passed as 32 bit input in 2's complement form
  reg clk;                  // sent clock pulse
  reg [10:0] i=0;           // the sample number is sent as an 11 bit binary value
  CLT abcd(.clk(clk), .Yin(Yin), .out(out), .i(i));     // instantiating the module CLT
    always #100 clk <= ~clk;
    initial begin 
        clk <= 0;
        #10 Yin =-32'd22; i= 11'd0;         /// yin has the input which is sent and i the sample number
        #200 Yin =-32'd18; i= 11'd1;
        #200 Yin =-32'd16; i= 11'd2;
        #200 Yin =-32'd14; i= 11'd3;
        #200 Yin =-32'd12; i= 11'd4;        // we have taken an actual ECG sample of 500 values and written C code
        #200 Yin =-32'd10; i= 11'd5;        // to generate this input of 500 samples in this format
        #200 Yin =-32'd8; i= 11'd6;
        #200 Yin =-32'd5; i= 11'd7;
        #200 Yin =-32'd2; i= 11'd8;
        #200 Yin =-32'd1; i= 11'd9;        // each sample has a delay of 200 units to provide sufficient calculation time
        #200 Yin =-32'd1; i= 11'd10;
        #200 Yin =-32'd2; i= 11'd11;
        #200 Yin =-32'd3; i= 11'd12;
        #200 Yin =-32'd3; i= 11'd13;
        #200 Yin =-32'd3; i= 11'd14;
        #200 Yin =-32'd2; i= 11'd15;
        #200 Yin =-32'd0; i= 11'd16;
        #200 Yin =32'd1; i= 11'd17;
        #200 Yin =32'd2; i= 11'd18;
        #200 Yin =32'd2; i= 11'd19;
        #200 Yin =32'd2; i= 11'd20;
        #200 Yin =32'd2; i= 11'd21;
        #200 Yin =32'd2; i= 11'd22;
        #200 Yin =32'd2; i= 11'd23;
        #200 Yin =32'd2; i= 11'd24;
        #200 Yin =32'd1; i= 11'd25;
        #200 Yin =32'd1; i= 11'd26;
        #200 Yin =32'd1; i= 11'd27;
        #200 Yin =32'd0; i= 11'd28;
        #200 Yin =32'd0; i= 11'd29;
        #200 Yin =32'd0; i= 11'd30;
        #200 Yin =32'd0; i= 11'd31;
        #200 Yin =32'd1; i= 11'd32;
        #200 Yin =32'd1; i= 11'd33;
        #200 Yin =32'd1; i= 11'd34;
        #200 Yin =32'd1; i= 11'd35;
        #200 Yin =32'd1; i= 11'd36;
        #200 Yin =32'd1; i= 11'd37;
        #200 Yin =32'd1; i= 11'd38;
        #200 Yin =32'd1; i= 11'd39;
        #200 Yin =32'd2; i= 11'd40;
        #200 Yin =32'd2; i= 11'd41;
        #200 Yin =32'd3; i= 11'd42;
        #200 Yin =32'd3; i= 11'd43;
        #200 Yin =32'd3; i= 11'd44;
        #200 Yin =32'd2; i= 11'd45;
        #200 Yin =32'd2; i= 11'd46;
        #200 Yin =32'd1; i= 11'd47;
        #200 Yin =32'd1; i= 11'd48;
        #200 Yin =32'd2; i= 11'd49;
        #200 Yin =32'd3; i= 11'd50;
        #200 Yin =32'd4; i= 11'd51;
        #200 Yin =32'd5; i= 11'd52;
        #200 Yin =32'd5; i= 11'd53;
        #200 Yin =32'd5; i= 11'd54;
        #200 Yin =32'd6; i= 11'd55;
        #200 Yin =32'd6; i= 11'd56;
        #200 Yin =32'd6; i= 11'd57;
        #200 Yin =32'd7; i= 11'd58;
        #200 Yin =32'd7; i= 11'd59;
        #200 Yin =32'd6; i= 11'd60;
        #200 Yin =32'd5; i= 11'd61;
        #200 Yin =32'd3; i= 11'd62;
        #200 Yin =32'd2; i= 11'd63;
        #200 Yin =32'd2; i= 11'd64;
        #200 Yin =32'd3; i= 11'd65;
        #200 Yin =32'd4; i= 11'd66;
        #200 Yin =32'd5; i= 11'd67;
        #200 Yin =32'd6; i= 11'd68;
        #200 Yin =32'd6; i= 11'd69;
        #200 Yin =32'd6; i= 11'd70;
        #200 Yin =32'd7; i= 11'd71;
        #200 Yin =32'd8; i= 11'd72;
        #200 Yin =32'd9; i= 11'd73;
        #200 Yin =32'd9; i= 11'd74;
        #200 Yin =32'd9; i= 11'd75;
        #200 Yin =32'd8; i= 11'd76;
        #200 Yin =32'd7; i= 11'd77;
        #200 Yin =32'd6; i= 11'd78;
        #200 Yin =32'd6; i= 11'd79;
        #200 Yin =32'd5; i= 11'd80;
        #200 Yin =32'd5; i= 11'd81;
        #200 Yin =32'd5; i= 11'd82;
        #200 Yin =32'd5; i= 11'd83;
        #200 Yin =32'd6; i= 11'd84;
        #200 Yin =32'd7; i= 11'd85;
        #200 Yin =32'd8; i= 11'd86;
        #200 Yin =32'd6; i= 11'd87;
        #200 Yin =32'd2; i= 11'd88;
        #200 Yin =-32'd4; i= 11'd89;
        #200 Yin =-32'd11; i= 11'd90;
        #200 Yin =-32'd15; i= 11'd91;
        #200 Yin =-32'd14; i= 11'd92;
        #200 Yin =-32'd9; i= 11'd93;
        #200 Yin =-32'd0; i= 11'd94;
        #200 Yin =32'd7; i= 11'd95;
        #200 Yin =32'd13; i= 11'd96;
        #200 Yin =32'd14; i= 11'd97;
        #200 Yin =32'd14; i= 11'd98;
        #200 Yin =32'd12; i= 11'd99;
        #200 Yin =32'd11; i= 11'd100;
        #200 Yin =32'd11; i= 11'd101;
        #200 Yin =32'd12; i= 11'd102;
        #200 Yin =32'd14; i= 11'd103;
        #200 Yin =32'd15; i= 11'd104;
        #200 Yin =32'd15; i= 11'd105;
        #200 Yin =32'd14; i= 11'd106;
        #200 Yin =32'd14; i= 11'd107;
        #200 Yin =32'd13; i= 11'd108;
        #200 Yin =32'd13; i= 11'd109;
        #200 Yin =32'd12; i= 11'd110;
        #200 Yin =32'd11; i= 11'd111;
        #200 Yin =32'd9; i= 11'd112;
        #200 Yin =32'd8; i= 11'd113;
        #200 Yin =32'd7; i= 11'd114;
        #200 Yin =32'd6; i= 11'd115;
        #200 Yin =32'd7; i= 11'd116;
        #200 Yin =32'd7; i= 11'd117;
        #200 Yin =32'd8; i= 11'd118;
        #200 Yin =32'd9; i= 11'd119;
        #200 Yin =32'd10; i= 11'd120;
        #200 Yin =32'd9; i= 11'd121;
        #200 Yin =32'd9; i= 11'd122;
        #200 Yin =32'd8; i= 11'd123;
        #200 Yin =32'd8; i= 11'd124;
        #200 Yin =32'd8; i= 11'd125;
        #200 Yin =32'd9; i= 11'd126;
        #200 Yin =32'd9; i= 11'd127;
        #200 Yin =32'd10; i= 11'd128;
        #200 Yin =32'd9; i= 11'd129;
        #200 Yin =32'd9; i= 11'd130;
        #200 Yin =32'd8; i= 11'd131;
        #200 Yin =32'd7; i= 11'd132;
        #200 Yin =32'd6; i= 11'd133;
        #200 Yin =32'd6; i= 11'd134;
        #200 Yin =32'd5; i= 11'd135;
        #200 Yin =32'd5; i= 11'd136;
        #200 Yin =32'd4; i= 11'd137;
        #200 Yin =32'd4; i= 11'd138;
        #200 Yin =32'd4; i= 11'd139;
        #200 Yin =32'd4; i= 11'd140;
        #200 Yin =32'd5; i= 11'd141;
        #200 Yin =32'd5; i= 11'd142;
        #200 Yin =32'd5; i= 11'd143;
        #200 Yin =32'd5; i= 11'd144;
        #200 Yin =32'd6; i= 11'd145;
        #200 Yin =32'd6; i= 11'd146;
        #200 Yin =32'd7; i= 11'd147;
        #200 Yin =32'd9; i= 11'd148;
        #200 Yin =32'd9; i= 11'd149;
        #200 Yin =32'd10; i= 11'd150;
        #200 Yin =32'd9; i= 11'd151;
        #200 Yin =32'd8; i= 11'd152;
        #200 Yin =32'd6; i= 11'd153;
        #200 Yin =32'd5; i= 11'd154;
        #200 Yin =32'd5; i= 11'd155;
        #200 Yin =32'd5; i= 11'd156;
        #200 Yin =32'd5; i= 11'd157;
        #200 Yin =32'd5; i= 11'd158;
        #200 Yin =32'd5; i= 11'd159;
        #200 Yin =32'd5; i= 11'd160;
        #200 Yin =32'd6; i= 11'd161;
        #200 Yin =32'd7; i= 11'd162;
        #200 Yin =32'd8; i= 11'd163;
        #200 Yin =32'd8; i= 11'd164;
        #200 Yin =32'd9; i= 11'd165;
        #200 Yin =32'd9; i= 11'd166;
        #200 Yin =32'd9; i= 11'd167;
        #200 Yin =32'd9; i= 11'd168;
        #200 Yin =32'd9; i= 11'd169;
        #200 Yin =32'd9; i= 11'd170;
        #200 Yin =32'd8; i= 11'd171;
        #200 Yin =32'd7; i= 11'd172;
        #200 Yin =32'd7; i= 11'd173;
        #200 Yin =32'd7; i= 11'd174;
        #200 Yin =32'd8; i= 11'd175;
        #200 Yin =32'd9; i= 11'd176;
        #200 Yin =32'd11; i= 11'd177;
        #200 Yin =32'd11; i= 11'd178;
        #200 Yin =32'd11; i= 11'd179;
        #200 Yin =32'd10; i= 11'd180;
        #200 Yin =32'd9; i= 11'd181;
        #200 Yin =32'd8; i= 11'd182;
        #200 Yin =32'd9; i= 11'd183;
        #200 Yin =32'd9; i= 11'd184;
        #200 Yin =32'd10; i= 11'd185;
        #200 Yin =32'd12; i= 11'd186;
        #200 Yin =32'd12; i= 11'd187;
        #200 Yin =32'd13; i= 11'd188;
        #200 Yin =32'd13; i= 11'd189;
        #200 Yin =32'd13; i= 11'd190;
        #200 Yin =32'd12; i= 11'd191;
        #200 Yin =32'd12; i= 11'd192;
        #200 Yin =32'd11; i= 11'd193;
        #200 Yin =32'd10; i= 11'd194;
        #200 Yin =32'd9; i= 11'd195;
        #200 Yin =32'd8; i= 11'd196;
        #200 Yin =32'd8; i= 11'd197;
        #200 Yin =32'd8; i= 11'd198;
        #200 Yin =32'd9; i= 11'd199;
        #200 Yin =32'd10; i= 11'd200;
        #200 Yin =32'd12; i= 11'd201;
        #200 Yin =32'd12; i= 11'd202;
        #200 Yin =32'd13; i= 11'd203;
        #200 Yin =32'd12; i= 11'd204;
        #200 Yin =32'd10; i= 11'd205;
        #200 Yin =32'd9; i= 11'd206;
        #200 Yin =32'd8; i= 11'd207;
        #200 Yin =32'd8; i= 11'd208;
        #200 Yin =32'd9; i= 11'd209;
        #200 Yin =32'd10; i= 11'd210;
        #200 Yin =32'd12; i= 11'd211;
        #200 Yin =32'd14; i= 11'd212;
        #200 Yin =32'd16; i= 11'd213;
        #200 Yin =32'd18; i= 11'd214;
        #200 Yin =32'd19; i= 11'd215;
        #200 Yin =32'd20; i= 11'd216;
        #200 Yin =32'd20; i= 11'd217;
        #200 Yin =32'd20; i= 11'd218;
        #200 Yin =32'd19; i= 11'd219;
        #200 Yin =32'd18; i= 11'd220;
        #200 Yin =32'd17; i= 11'd221;
        #200 Yin =32'd17; i= 11'd222;
        #200 Yin =32'd17; i= 11'd223;
        #200 Yin =32'd17; i= 11'd224;
        #200 Yin =32'd16; i= 11'd225;
        #200 Yin =32'd15; i= 11'd226;
        #200 Yin =32'd14; i= 11'd227;
        #200 Yin =32'd12; i= 11'd228;
        #200 Yin =32'd12; i= 11'd229;
        #200 Yin =32'd12; i= 11'd230;
        #200 Yin =32'd12; i= 11'd231;
        #200 Yin =32'd13; i= 11'd232;
        #200 Yin =32'd12; i= 11'd233;
        #200 Yin =32'd11; i= 11'd234;
        #200 Yin =32'd10; i= 11'd235;
        #200 Yin =32'd9; i= 11'd236;
        #200 Yin =32'd8; i= 11'd237;
        #200 Yin =32'd9; i= 11'd238;
        #200 Yin =32'd10; i= 11'd239;
        #200 Yin =32'd12; i= 11'd240;
        #200 Yin =32'd12; i= 11'd241;
        #200 Yin =32'd12; i= 11'd242;
        #200 Yin =32'd11; i= 11'd243;
        #200 Yin =32'd10; i= 11'd244;
        #200 Yin =32'd9; i= 11'd245;
        #200 Yin =32'd8; i= 11'd246;
        #200 Yin =32'd8; i= 11'd247;
        #200 Yin =32'd8; i= 11'd248;
        #200 Yin =32'd8; i= 11'd249;
        #200 Yin =32'd8; i= 11'd250;
        #200 Yin =32'd7; i= 11'd251;
        #200 Yin =32'd5; i= 11'd252;
        #200 Yin =32'd4; i= 11'd253;
        #200 Yin =32'd3; i= 11'd254;
        #200 Yin =32'd3; i= 11'd255;
        #200 Yin =32'd4; i= 11'd256;
        #200 Yin =32'd4; i= 11'd257;
        #200 Yin =32'd4; i= 11'd258;
        #200 Yin =32'd3; i= 11'd259;
        #200 Yin =32'd1; i= 11'd260;
        #200 Yin =32'd0; i= 11'd261;
        #200 Yin =-32'd0; i= 11'd262;
        #200 Yin =-32'd0; i= 11'd263;
        #200 Yin =-32'd0; i= 11'd264;
        #200 Yin =-32'd0; i= 11'd265;
        #200 Yin =-32'd0; i= 11'd266;
        #200 Yin =-32'd0; i= 11'd267;
        #200 Yin =-32'd1; i= 11'd268;
        #200 Yin =-32'd1; i= 11'd269;
        #200 Yin =-32'd1; i= 11'd270;
        #200 Yin =-32'd1; i= 11'd271;
        #200 Yin =-32'd1; i= 11'd272;
        #200 Yin =-32'd1; i= 11'd273;
        #200 Yin =-32'd1; i= 11'd274;
        #200 Yin =-32'd1; i= 11'd275;
        #200 Yin =-32'd0; i= 11'd276;
        #200 Yin =-32'd0; i= 11'd277;
        #200 Yin =32'd0; i= 11'd278;
        #200 Yin =32'd0; i= 11'd279;
        #200 Yin =32'd1; i= 11'd280;
        #200 Yin =32'd1; i= 11'd281;
        #200 Yin =32'd1; i= 11'd282;
        #200 Yin =32'd0; i= 11'd283;
        #200 Yin =-32'd0; i= 11'd284;
        #200 Yin =-32'd1; i= 11'd285;
        #200 Yin =-32'd1; i= 11'd286;
        #200 Yin =-32'd0; i= 11'd287;
        #200 Yin =32'd0; i= 11'd288;
        #200 Yin =32'd0; i= 11'd289;
        #200 Yin =32'd1; i= 11'd290;
        #200 Yin =32'd0; i= 11'd291;
        #200 Yin =-32'd0; i= 11'd292;
        #200 Yin =-32'd0; i= 11'd293;
        #200 Yin =-32'd0; i= 11'd294;
        #200 Yin =32'd0; i= 11'd295;
        #200 Yin =32'd1; i= 11'd296;
        #200 Yin =32'd1; i= 11'd297;
        #200 Yin =32'd0; i= 11'd298;
        #200 Yin =-32'd1; i= 11'd299;
        #200 Yin =-32'd3; i= 11'd300;
        #200 Yin =-32'd5; i= 11'd301;
        #200 Yin =-32'd6; i= 11'd302;
        #200 Yin =-32'd6; i= 11'd303;
        #200 Yin =-32'd5; i= 11'd304;
        #200 Yin =-32'd4; i= 11'd305;
        #200 Yin =-32'd3; i= 11'd306;
        #200 Yin =-32'd1; i= 11'd307;
        #200 Yin =32'd0; i= 11'd308;
        #200 Yin =32'd2; i= 11'd309;
        #200 Yin =32'd5; i= 11'd310;
        #200 Yin =32'd7; i= 11'd311;
        #200 Yin =32'd9; i= 11'd312;
        #200 Yin =32'd10; i= 11'd313;
        #200 Yin =32'd12; i= 11'd314;
        #200 Yin =32'd13; i= 11'd315;
        #200 Yin =32'd16; i= 11'd316;
        #200 Yin =32'd19; i= 11'd317;
        #200 Yin =32'd22; i= 11'd318;
        #200 Yin =32'd23; i= 11'd319;
        #200 Yin =32'd21; i= 11'd320;
        #200 Yin =32'd18; i= 11'd321;
        #200 Yin =32'd13; i= 11'd322;
        #200 Yin =32'd9; i= 11'd323;
        #200 Yin =32'd6; i= 11'd324;
        #200 Yin =32'd5; i= 11'd325;
        #200 Yin =32'd6; i= 11'd326;
        #200 Yin =32'd8; i= 11'd327;
        #200 Yin =32'd10; i= 11'd328;
        #200 Yin =32'd10; i= 11'd329;
        #200 Yin =32'd8; i= 11'd330;
        #200 Yin =32'd4; i= 11'd331;
        #200 Yin =-32'd1; i= 11'd332;
        #200 Yin =-32'd9; i= 11'd333;
        #200 Yin =-32'd19; i= 11'd334;
        #200 Yin =-32'd28; i= 11'd335;
        #200 Yin =-32'd35; i= 11'd336;
        #200 Yin =-32'd36; i= 11'd337;
        #200 Yin =-32'd33; i= 11'd338;
        #200 Yin =-32'd25; i= 11'd339;
        #200 Yin =-32'd15; i= 11'd340;
        #200 Yin =-32'd5; i= 11'd341;
        #200 Yin =32'd1; i= 11'd342;
        #200 Yin =32'd4; i= 11'd343;
        #200 Yin =32'd5; i= 11'd344;
        #200 Yin =32'd5; i= 11'd345;
        #200 Yin =32'd4; i= 11'd346;
        #200 Yin =32'd3; i= 11'd347;
        #200 Yin =32'd3; i= 11'd348;
        #200 Yin =32'd4; i= 11'd349;
        #200 Yin =32'd4; i= 11'd350;
        #200 Yin =32'd5; i= 11'd351;
        #200 Yin =32'd5; i= 11'd352;
        #200 Yin =32'd4; i= 11'd353;
        #200 Yin =32'd2; i= 11'd354;
        #200 Yin =32'd0; i= 11'd355;
        #200 Yin =-32'd1; i= 11'd356;
        #200 Yin =-32'd3; i= 11'd357;
        #200 Yin =-32'd3; i= 11'd358;
        #200 Yin =-32'd2; i= 11'd359;
        #200 Yin =-32'd0; i= 11'd360;
        #200 Yin =32'd1; i= 11'd361;
        #200 Yin =32'd3; i= 11'd362;
        #200 Yin =32'd3; i= 11'd363;
        #200 Yin =32'd2; i= 11'd364;
        #200 Yin =32'd0; i= 11'd365;
        #200 Yin =-32'd1; i= 11'd366;
        #200 Yin =-32'd1; i= 11'd367;
        #200 Yin =-32'd2; i= 11'd368;
        #200 Yin =-32'd1; i= 11'd369;
        #200 Yin =-32'd1; i= 11'd370;
        #200 Yin =-32'd1; i= 11'd371;
        #200 Yin =-32'd2; i= 11'd372;
        #200 Yin =-32'd3; i= 11'd373;
        #200 Yin =-32'd4; i= 11'd374;
        #200 Yin =-32'd5; i= 11'd375;
        #200 Yin =-32'd4; i= 11'd376;
        #200 Yin =-32'd3; i= 11'd377;
        #200 Yin =-32'd3; i= 11'd378;
        #200 Yin =-32'd2; i= 11'd379;
        #200 Yin =-32'd2; i= 11'd380;
        #200 Yin =-32'd2; i= 11'd381;
        #200 Yin =-32'd2; i= 11'd382;
        #200 Yin =-32'd1; i= 11'd383;
        #200 Yin =-32'd1; i= 11'd384;
        #200 Yin =-32'd0; i= 11'd385;
        #200 Yin =-32'd1; i= 11'd386;
        #200 Yin =-32'd1; i= 11'd387;
        #200 Yin =-32'd1; i= 11'd388;
        #200 Yin =-32'd2; i= 11'd389;
        #200 Yin =-32'd2; i= 11'd390;
        #200 Yin =-32'd3; i= 11'd391;
        #200 Yin =-32'd3; i= 11'd392;
        #200 Yin =-32'd4; i= 11'd393;
        #200 Yin =-32'd4; i= 11'd394;
        #200 Yin =-32'd5; i= 11'd395;
        #200 Yin =-32'd5; i= 11'd396;
        #200 Yin =-32'd6; i= 11'd397;
        #200 Yin =-32'd6; i= 11'd398;
        #200 Yin =-32'd6; i= 11'd399;
        #200 Yin =-32'd6; i= 11'd400;
        #200 Yin =-32'd5; i= 11'd401;
        #200 Yin =-32'd4; i= 11'd402;
        #200 Yin =-32'd3; i= 11'd403;
        #200 Yin =-32'd2; i= 11'd404;
        #200 Yin =-32'd1; i= 11'd405;
        #200 Yin =-32'd0; i= 11'd406;
        #200 Yin =-32'd1; i= 11'd407;
        #200 Yin =-32'd1; i= 11'd408;
        #200 Yin =-32'd2; i= 11'd409;
        #200 Yin =-32'd3; i= 11'd410;
        #200 Yin =-32'd4; i= 11'd411;
        #200 Yin =-32'd4; i= 11'd412;
        #200 Yin =-32'd4; i= 11'd413;
        #200 Yin =-32'd4; i= 11'd414;
        #200 Yin =-32'd3; i= 11'd415;
        #200 Yin =-32'd3; i= 11'd416;
        #200 Yin =-32'd2; i= 11'd417;
        #200 Yin =-32'd2; i= 11'd418;
        #200 Yin =-32'd2; i= 11'd419;
        #200 Yin =-32'd2; i= 11'd420;
        #200 Yin =-32'd1; i= 11'd421;
        #200 Yin =-32'd1; i= 11'd422;
        #200 Yin =-32'd1; i= 11'd423;
        #200 Yin =-32'd1; i= 11'd424;
        #200 Yin =-32'd2; i= 11'd425;
        #200 Yin =-32'd2; i= 11'd426;
        #200 Yin =-32'd3; i= 11'd427;
        #200 Yin =-32'd2; i= 11'd428;
        #200 Yin =-32'd2; i= 11'd429;
        #200 Yin =-32'd1; i= 11'd430;
        #200 Yin =-32'd0; i= 11'd431;
        #200 Yin =-32'd0; i= 11'd432;
        #200 Yin =-32'd0; i= 11'd433;
        #200 Yin =-32'd1; i= 11'd434;
        #200 Yin =-32'd1; i= 11'd435;
        #200 Yin =-32'd1; i= 11'd436;
        #200 Yin =-32'd0; i= 11'd437;
        #200 Yin =32'd0; i= 11'd438;
        #200 Yin =32'd0; i= 11'd439;
        #200 Yin =32'd1; i= 11'd440;
        #200 Yin =32'd1; i= 11'd441;
        #200 Yin =32'd1; i= 11'd442;
        #200 Yin =32'd0; i= 11'd443;
        #200 Yin =32'd0; i= 11'd444;
        #200 Yin =-32'd0; i= 11'd445;
        #200 Yin =-32'd0; i= 11'd446;
        #200 Yin =-32'd0; i= 11'd447;
        #200 Yin =-32'd1; i= 11'd448;
        #200 Yin =-32'd1; i= 11'd449;
        #200 Yin =-32'd1; i= 11'd450;
        #200 Yin =-32'd1; i= 11'd451;
        #200 Yin =-32'd1; i= 11'd452;
        #200 Yin =-32'd1; i= 11'd453;
        #200 Yin =-32'd1; i= 11'd454;
        #200 Yin =-32'd1; i= 11'd455;
        #200 Yin =-32'd0; i= 11'd456;
        #200 Yin =32'd0; i= 11'd457;
        #200 Yin =32'd0; i= 11'd458;
        #200 Yin =32'd0; i= 11'd459;
        #200 Yin =32'd0; i= 11'd460;
        #200 Yin =-32'd0; i= 11'd461;
        #200 Yin =-32'd0; i= 11'd462;
        #200 Yin =-32'd1; i= 11'd463;
        #200 Yin =-32'd1; i= 11'd464;
        #200 Yin =-32'd2; i= 11'd465;
        #200 Yin =-32'd3; i= 11'd466;
        #200 Yin =-32'd4; i= 11'd467;
        #200 Yin =-32'd4; i= 11'd468;
        #200 Yin =-32'd3; i= 11'd469;
        #200 Yin =-32'd2; i= 11'd470;
        #200 Yin =-32'd0; i= 11'd471;
        #200 Yin =32'd2; i= 11'd472;
        #200 Yin =32'd4; i= 11'd473;
        #200 Yin =32'd6; i= 11'd474;
        #200 Yin =32'd7; i= 11'd475;
        #200 Yin =32'd7; i= 11'd476;
        #200 Yin =32'd7; i= 11'd477;
        #200 Yin =32'd7; i= 11'd478;
        #200 Yin =32'd6; i= 11'd479;
        #200 Yin =32'd4; i= 11'd480;
        #200 Yin =32'd3; i= 11'd481;
        #200 Yin =32'd1; i= 11'd482;
        #200 Yin =32'd0; i= 11'd483;
        #200 Yin =32'd0; i= 11'd484;
        #200 Yin =-32'd0; i= 11'd485;
        #200 Yin =32'd0; i= 11'd486;
        #200 Yin =32'd0; i= 11'd487;
        #200 Yin =32'd1; i= 11'd488;
        #200 Yin =32'd3; i= 11'd489;
        #200 Yin =32'd5; i= 11'd490;
        #200 Yin =32'd7; i= 11'd491;
        #200 Yin =32'd0; i= 11'd492;
        #200 Yin =32'd0; i= 11'd493;
        #200 Yin =32'd0; i= 11'd494;
        #200 Yin =32'd0; i= 11'd495;
        #200 Yin =32'd0; i= 11'd496;
        #200 Yin =32'd0; i= 11'd497;
        #200 Yin =32'd0; i= 11'd498;
        #200 Yin =32'd0; i= 11'd499;
        #200 Yin =-32'd0; i= 11'd500;
    end
endmodule